`ifndef ALU_MATRIX_DEFINES
`define ALU_MATRIX_DEFINES


`define AXI_DATA_W   8
`define APB_ADDR_W   32
`define APB_DATA_W   32
`define BUFFER_DEPTH 64

`define MAX_DET_RANK 8

`endif // !ALU_MATRIX_DEFINES