`ifndef IRQ_AGENT_IF
`define IRQ_AGENT_IF

interface irq_agent_if();

  logic irq;
  
endinterface

`endif //!IRQ_AGENT_IF
